//регситр результата (сдвиговый + очистка)
module rr (data, load, en, clk, r, rr_out); 	//объявление модуля и его входов/выходов
	parameter N = 4;									//параметр для изменения размера шины данных
	input wire [(2*N-1):0] data;					//вход - шина 2N
   input load; 										//разрешение записи
	input en;											//разрешение
	input clk;											//тактовый сигнал
	input r;												//сброс
	output reg [(2*N-1):0] rr_out; 				//выход - 2N

	reg [(2*N-1):0] state;							//внутренний регистр состояния
	
	always @ (posedge clk)							//блок описания поведения, чувствительный к изменению сигнала clk по положительому фронту (posedge)
	begin
		if (r) begin									//если r = 1
			state = 0;									//сброс в 0
			end
		else if (en) begin							//если есть разрешение
			if (load) begin							//если разрешена запись
				state = data;							//запись входящих данных
				end		
			else begin									//иначе (сдвиг)
				state = {state[2*N-2:0], state[2*N-1]};	//сдвиг на 1 бил влево, младший бит принимает значение знакового бита
			end
		end
		rr_out = state;								//передача state на выход регистра (без условий, каждый раз при изменении clk по положительному фронту)
	end
endmodule 
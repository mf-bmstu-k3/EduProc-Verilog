//кс2 - формирование признака результата
module ks3 (rr, ks3_out);					//объявление модуля и его входов/выходов
	parameter N = 4;							//параметр для изменения размера шины данных
	input wire [N:0] rr;   					//вход данных с регистра результата
	output reg [1:0] ks3_out;   			//регистр данных (2 бита) - выход
	
	wire [(2*N):0] zero = 0;				//2N-битный 0
	
	always @* begin							//блок описания поведения комбинационной схемы
		ks3_out[0] = rr[4]|(rr[3]);
		ks3_out[1] = {((~rr[4]|(~rr[3]))&(rr[4]|rr[3]|rr[2]|rr[1]|rr[0]))};
	end

endmodule 


module BO_as_one_module (clk, a, b, y, rr, priznak, f);
	parameter N = 4; //параметр, задает разрядность операндов
	
	input clk;								//тактовый сигнал
	input wire [(N-1):0] a; 			//первый операнд
	input wire [(N-1):0] b; 			//второй операнд
	input wire [10:1] y; 				//управляющие сигналы
	output reg [(2*N-1):0] rr; 		//результат
	output reg [1:0] priznak; 			//признак результата
	output reg [2:0] f; 					//признак отрицательного нуля, анализируемый разряд множителя, знак множителя

												//внутрение регистры
	reg [(N-1):0] RA; 					//а
	reg [(N-1):0] RB; 					//в
	reg [(2*N):0] zero = 0; 			//0 (вспомогательный)
												
												//комбинационные схемы
	reg [(2*N-1):0] d; 					//выход КС1
	reg [(2*N-1):0] q; 					//выход КС2
	reg [(2*N-1):0] s; 					//выход сумматора
	reg [1:0] pr; 							//выход КС3

				
	//этот процесс описывает логику работы регистра RA 
	always @(posedge clk) begin		//по положительному фронту clk
		if (y[1]) begin 					//если есть разрешение
			RA = a;							//выполняется прием первого операнда
		end
	end
	
	//этот процесс описывает логику работы регистра RB 
	always @(posedge clk) begin		//по положительному фронту clk
		if (y[3]) begin 					//если есть разрешение тактирования
			if (y[2]) begin				//если разрешена загрузка
				RB = b;  					//прием второго операнда
			end
			else begin
				RB = {RB[N-1], RB[(N-3):0], 1'b0}; //иначе сдвиг влево RB с сохранением знака
			end
		end
	end
	
	//этот процесс описывает КС1
	//d - выход КС1
	always @* begin
		case (y[5:4])
			2'b01: begin 										//если y4=1
				if (RA[N-1]) begin							//если число отрицательное
					d[(2*N-1):N] = ~zero[(2*N-1):N];		//старшим разрядам присваивается 1
				end
				else if (!RA[N-1]) begin					//иначе если число положительное
					d[(2*N-1):N] = zero[(2*N-1):N];		//старшим разрядам присваивается 0
				end
				d[(N-1):0] = RA;								//передаем на суммирование +А
			end
			2'b10: begin
				if (RA[N-1]) begin							//если число отрицательное
					d[(2*N-1):N] = zero[(2*N-1):N];		//старшим разрядам присваивается0
				end
				else if (!RA[N-1]) begin					//иначе если число положительное
					d[(2*N-1):N] = ~zero[(2*N-1):N];		//старшим разрядам присваивается 1
				end
				d[(N-1):0] = ~RA;								//передаем на суммирование -А
			end
			default: begin
				d[(2*N-1):0] = 0;		//ноль в остальных случаях
			end
		endcase
	end
	
	//этот процесс описывает КС2
	//q - выход КС2
	always @* begin
		if(y[9]) begin
				q[(2*N-1):0] = rr[(2*N-1):0];
		end
		else begin
			if (RB[N-1]) begin							
				q[(2*N-1):N] = ~zero[(2*N-1):N];		
			end
			else if (!RB[N-1]) begin					
				q[(2*N-1):N] = zero[(2*N-1):N];		
			end
			q[(N-1):0] = RB[(N-1):0];		
		end
	end
	
	
	//этот процесс описывает работу сумматора в обратном коде
	//к его входам подключены выходы КС1 и КС2
	reg [(2*N):0] sym = 0; 	//для вычисления суммы
	
	always @* begin
		sym = d + q;			//сложение
		sym[(2*N-1):0] = sym + sym[2*N];
		s <= sym[(2*N-1):0];
	end
	
	//этот процесс описывает работу регистра результата
	always @(posedge clk) begin
		if (y[8]) begin
			rr = zero;   				//очистка rr
		end
		else if (y[7]) begin 		//если есть разрешение тактирования
			if (y[6]) begin 
				rr = s;					//загрузка rr
			end
			else begin
				rr = {rr[(2*N-2):0], rr[2*N-1]}; //циклический сдвиг влево rr
			end
		end
	end
	
	//этот процесс описывает КС3, которая формирует признак результата
	//q - выход КС2
	always @* begin
		pr[0] = rr[4]|(rr[3]);
		pr[1] = {((~rr[4]|(~rr[3]))&(rr[4]|rr[3]|rr[2]|rr[1]|rr[0]))};
	end

	//этот процесс описывает работу регистра признака
	always @(posedge clk) begin
		if (y[10]) begin 
			priznak<=pr; 							//запоминаем признак результата
		end
	end
	
	//ниже приводится описание логических условий
	always @* begin
		f[0]= RB[N-1];   							//знак множителя
		f[1]= RB[N-2];								//анализируемый разряд множителя
		if (rr[N:0]==(~zero[N:0])) begin		//отрицательный ноль
			f[2]= 1'b1;
		end
		else begin
			f[2]= 1'b0;			
		end
	end
	
endmodule
//сдвиговый регистр (б)
module rb (data, load, clk, en, rb_out); 				//объявление модуля и его входов/выходов
	parameter N = 4;											//параметр для изменения размера шины данных
	input wire [(N-1):0] data;								//шина входящих данных
	input load;													//разрешение записи
   input clk; 													//тактовый сигнал
	input en;													//разрешение
	output reg [(N-1):0] rb_out;  						//регистр данных (выход)

	reg [(N-1):0] state;										//внутренний регистр данных
	
	always @ (posedge clk)									//блок описания поведения, чувствительный к изменению сигнала clk по положительому фронту (posedge)
	begin												
		if (en) begin											//если en = 1
			if (load) begin									//если load = 1 (запись разрешена)
				state = data;									//state принимает значение data 
			end
			else if (!load) begin							//если load = 0 (запись запрещена = сдвиг)
				state = {state[N-1], state[(N-3):0], 1'b0}; 	//сдвиг регистра влево с сохранением знакового разряда
																	//конструкцией state = {a, b, c} мы задаем каждый бит шины по очереди, начиная со старших битов
																	// было	state [N] 	state [N-1] ..... state [1] state [0]
																	//стало	state [N-1]	state [N-2] ..... state [0]    0
			end
		end
		rb_out = state;										//передача state на выход регистра (без условий, каждый раз при изменении clk по положительному фронту)
	end
endmodule 



//регистр признака результата (аналогичен регстру а, но имеет фиксированный размер)
module rpr (data, clk, en, ra_out);	//объявление модуля и его входов/выходов
	input wire [1:0] data;				//вход - два бита данных
   input clk;								//тактовый сигнал
	input en;								//разрешенеие
	output reg [1:0] ra_out;   		//выход - два бита данных
	
	always @*								//блок описания поведения комбинационной схемы
	begin
		if (en) begin						//если разрешение = 1
			ra_out = data;					//выход = вход
		end
	end
endmodule 
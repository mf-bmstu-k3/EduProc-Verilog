// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Mon Apr 22 11:28:20 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,x[2:0],sno,i[1:0],
    y[9:0],sko,incr_i);

    input reset;
    input clock;
    input [2:0] x;
    input sno;
    input [1:0] i;
    tri0 reset;
    tri0 [2:0] x;
    tri0 sno;
    tri0 [1:0] i;
    output [9:0] y;
    output sko;
    output incr_i;
    reg [9:0] y;
    reg sko;
    reg incr_i;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter s0=0,s1=1,s2=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or x or sno or i)
    begin
        if (reset) begin
            reg_fstate <= s0;
            y <= 10'b0000000000;
            sko <= 1'b0;
            incr_i <= 1'b0;
        end
        else begin
            y <= 10'b0000000000;
            sko <= 1'b0;
            incr_i <= 1'b0;
            case (fstate)
                s0: begin
                    if (~(sno))
                        reg_fstate <= s0;
                    else if (sno)
                        reg_fstate <= s1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s0;

                    sko <= 1'b0;

                    if (~(sno))
                        y <= 10'b0000000000;
                    else if (sno)
                        y <= 10'b0011000111;
                    // Inserting 'else' block to prevent latch inference
                    else
                        y <= 10'b0000000000;
                end
                s1: begin
                    reg_fstate <= s2;

                    sko <= 1'b0;

                    if ((x[1] & ~(x[0])))
                        y <= 10'b0001101000;
                    else if ((~(x[1]) & x[0]))
                        y <= 10'b0001110000;
                    else
                        y <= 10'b0001100000;
                end
                s2: begin
                    if ((i[1:0] == 2'b11))
                        reg_fstate <= s0;
                    else if ((i[1:0] != 2'b11))
                        reg_fstate <= s1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s2;

                    if ((i[1:0] == 2'b11))
                        sko <= 1'b1;
                    else if ((i[1:0] != 2'b11))
                        sko <= 1'b0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        sko <= 1'b0;

                    if ((i[1:0] != 2'b11))
                        incr_i <= 1'b1;
                    else
                        incr_i <= 1'b0;

                    if ((i[1:0] != 2'b11))
                        y <= 10'b0001000100;
                    else if ((i[1:0] == 2'b11))
                        y <= 10'b0000000000;
                    // Inserting 'else' block to prevent latch inference
                    else
                        y <= 10'b0000000000;
                end
                default: begin
                    y <= 10'bxxxxxxxxxx;
                    sko <= 1'bx;
                    incr_i <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1

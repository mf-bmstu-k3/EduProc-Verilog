//кс2 - передача на сумматор значение б или значение результата
module ks2 (rr, rb, y9, ks2_out);						//объявление модуля и его входов/выходов
	parameter N = 4;											//параметр для изменения размера шины данных
	input wire [(2*N-1):0] rr;   							//вход данных с регистра результата (2N бит)
	input wire [(N-1):0] rb; 								//вход данных с регистра б (N бит)
   input y9; 													//управляющий сигнал
	output reg [(2*N-1):0] ks2_out;   					//выход - регистр данных (2N бит)
	
	integer i;                                      //инкремент для счетчика
	
	always @* begin											//блок описания поведения комбинационной схемы
		if (y9 == 0) begin                          	//если y9 = 0 (сложение)
			for (i = 0; i < 2*N; i = i + 1) begin   	//цикл от 0 до 2N
				if (i < N) begin                    	
					ks2_out[i] = {rb[i]};           		//младшим разрядам присваивается значение RB
				end
				if (i >= N) begin	
					ks2_out[i] = {rb[N-1]};         		//старшим разрядам присваивается значение знакового бита RB
				end                          
			end
		end
		else begin                                  	//y9 = 1 - умножение
			for (i = 0; i < 2*N; i = i + 1) begin   	//цикл от 0 до 2N
				ks2_out[i] = {rr[i]};               	//передача регистра результатаЫ
				end
		end
	end
endmodule 
//сумматор
module sum (a, b, sum_out);			//объявление модуля и его входов/выходов
	parameter N = 4;						//параметр для изменения размера шины данных
	input unsigned [(2*N-1):0] a;		//вход данных с регистра А (2N)
	input unsigned [(2*N-1):0] b;		//вход данных с регистра Б (2N)
	output reg [(2*N-1):0] sum_out;	//выход (2N)
		
	reg [(2*N-1):0] sym;					//вгутренний регистр суммы
	reg carry;								//регистр для бита переноса
	
	always @*								//блок описания поведения комбинационной схемы
	begin
		{carry, sym} = a+b;				//запись суммы и бита переноса
		sum_out = sym + carry;			//вывод суммы с учетом переноса
	end
endmodule 




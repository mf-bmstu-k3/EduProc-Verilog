//кс1 - передача на сумматор +-РА
module ks1 (ra, y4, y5, ks1_out);						//объявление модуля и его входов/выходов
	parameter N = 4;											//параметр для изменения размера шины данных
	input wire [(N-1):0] ra;								//вход данных с ра (N бит)
   input y4;    												//управляющий сигналы
   input y5; 
	output reg [(2*N-1):0] ks1_out;   					//выход данных (2N бит)

	reg [(2*N-1):0] zero = 0; 								//регистр в котором хранится 2N-разрядный 0
																	//этот регистр нужен чтобы заполнять знаковым разрядом биты с 2N по N+1 /
																	//для заполнения 0м используется регистр без изменений, для 1 - инвертированный
																	
	always @*													//блок описания поведения комбинационной схемы
	begin
		if (y4) begin											//если включена передача +RA
			if (ra[N-1]) begin								//если число отрицательное
				ks1_out[(2*N-1):N] = ~zero[(2*N-1):N];	//старшим разрядам присваивается не 0, т.е. 1
			end
			else if (!ra[N-1]) begin						//иначе если число положительное
				ks1_out[(2*N-1):N] = zero[(2*N-1):N];	//старшим разрядам присваивается 0
			end
			ks1_out[(N-1):0] = ra[(N-1):0];				//младшим разрядам присваивается значение RA
		end
		else if (y5) begin									//если включена передача -RA
			if (ra[N-1]) begin								//если число отрицательное
				ks1_out[(2*N-1):N] = zero[(2*N-1):N];	//старшим разрядам присваивается 0
			end
			else if (!ra[N-1]) begin						//иначе если число положительное
				ks1_out[(2*N-1):N] = ~zero[(2*N-1):N]; //старшим разрядам присваивается 1
			end
			ks1_out[(N-1):0] = ~ra[(N-1):0];				//младшим разрядам присваивается не RA
		end
		else if (!(y4+y5)) begin							//если y4 и y5 равны нулю
			ks1_out = zero;									//0 на выходе
		end			
	end
endmodule 
//запоминающий регистр (а, результат)
module reg_r (data, clk, en, reg_out); 	//объявление модуля и его входов/выходов
	parameter N = 4;								//параметр для изменения размера шины данных
														//описание входов и выходов модуля
	input wire [(N-1):0] data;					//шина входящих данных (N бит)
   input clk;										//тактовый сигнал
	input en;										//разрешение записи
	output reg [(N-1):0] reg_out;   			//выход модуля, регистр на N бит
	
	always @ (posedge clk)						//блок описания поведения, чувствительный к изменению сигнала clk по положительому фронту (posedge)
	begin												
		if (en) begin								//если на разрешающем входе "1"
			reg_out <= data;						//регистру ra_out присваивается значение входа data
		end							
	end
	
endmodule 



